../tb/pat//my_seq.sv