../tb/pat/test_burst_transfer/my_seq.sv