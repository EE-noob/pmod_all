../tb/pat/test_burst_transfer/my_test.sv