../tb/pat/test_single_transfer/my_seq.sv