../tb/pat/test_single_transfer/my_test.sv