../tb/pat//my_test.sv