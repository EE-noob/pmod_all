../tb/pat/mult_wr_trans/my_seq.sv