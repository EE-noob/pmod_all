  `ifndef _AXI_UART_DEFINES_H_
  `define _AXI_UART_DEFINES_H_

  `define _AXI_UART_DATA_WIDTH_ 32
  `define _AXI_UART_ADDR_WIDTH_ 5
  `define _AXI_UART_FIFO_DEPTH_ 16//32
  `define _AXI_UART_DIV_WIDTH_  32
  `define _AXI_UART_RESP_WIDTH_ 2
  `define _AXI_UART_ID_WIDTH_   12

  `define _AXI_UART_DEADLOCK_   2**20

  `endif
